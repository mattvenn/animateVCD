localparam NOP         = 0; //1
localparam LD_DATA     = 1; //2
localparam LD_COEFF    = 2; //4
localparam ADD         = 3; //8
localparam MULT        = 4; //16
localparam WRITE       = 5; //32
