localparam NOP         = 0;
localparam MEM1        = 1;
localparam MEM2        = 2;
localparam ADD         = 3;
localparam MULT        = 4;
localparam WRITE       = 5;
